module Encoder_4to2(
	input  [3:0] in,
	output [1:0] out
);
/*
------------------------------------------------
   in[3]  in[2]  in[1]  in[0] | out[1] out[0]  
------------------------------------------------
    1      1      0      1    |   0      0  
    1      1      1      0    |   0      1  
    0      1      1      0    |   1      0   
	 0      0      0      1    |   1      1        

*/
 
assign out[0] = ~in[2] | (~in[0] & in[3]);
assign out[1] = ~in[3];

endmodule 